module sqrt64(
    input clk,
    input unsigned [63:0] in,
    output unsigned [31:0] out
);


endmodule
