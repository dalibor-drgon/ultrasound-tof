module atan2(
    input clk,
    input y_neg, y_zero,
    input [20:0] y_log,
    input x_neg, x_zero,
    input [20:0] x_log
);

    

endmodule
